`define WR_DATA_WIDTH_MUL 1 // WR_DATA_WIDTH = WR_DATA_WIDTH_MUL * DATA_WIDTH
`define RD_DATA_WIDTH_MUL 1 // RD_DATA_WIDTH = RD_DATA_WIDTH_MUL * DATA_WIDTH
`define DATA_WIDTH 8 
`define ADDRESS_WIDTH 4
`define WR_DATA_WIDTH `WR_DATA_WIDTH_MUL * `DATA_WIDTH
`define RD_DATA_WIDTH `RD_DATA_WIDTH_MUL * `DATA_WIDTH
`define FIFO_DEPTH (1 << `ADDRESS_WIDTH)
`define WR_COUNT 17
`define RD_COUNT 17
`define HALF_PERIOD_WRCLK 15
`define HALF_PERIOD_RDCLK 18